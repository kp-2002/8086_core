module exe_unit(
	);

	

endmodule
