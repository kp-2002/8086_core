module 8086_core_top(
	);



endmodule
