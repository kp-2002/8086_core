module bus_if_unit(
	
	);

	

endmodule	
